library verilog;
use verilog.vl_types.all;
entity tb_parteIII is
end tb_parteIII;
